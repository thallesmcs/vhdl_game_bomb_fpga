----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    19:51:11 06/14/2023 
-- Design Name: 
-- Module Name:    imp - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity imp is
    Port ( clock, btn3, btn1 : in  STD_LOGIC;
           switch : in  STD_LOGIC_VECTOR (7 downto 0);
           led : out  STD_LOGIC_VECTOR (7 downto 0);
           cx : out  STD_LOGIC_VECTOR (7 downto 0);
           an : out  STD_LOGIC_VECTOR (3 downto 0));
end imp;

architecture Behavioral of imp is

signal clk_1, clk_250, clk_3 : STD_LOGIC;

signal q_nc, qc, q_nr, qr, binario_aleatorio : STD_LOGIC_VECTOR(7 downto 0);
signal sw_s : STD_LOGIC_VECTOR(7 downto 0);
signal led_s : STD_LOGIC_VECTOR(7 downto 0);
signal an_s : STD_LOGIC_VECTOR(3 downto 0);
signal cx_s : STD_LOGIC_VECTOR(7 downto 0);
signal disp0, disp1, disp2, disp3 : STD_LOGIC_VECTOR(7 downto 0);
signal confirmador, btn_s: STD_LOGIC;
signal chave: STD_LOGIC := '1';

component div_f is
    Port (clk_d, reset : in STD_LOGIC;
			clk_1, clk_250, clk_3 : out STD_LOGIC);
end component;


component countdowni is
	port(clock : in STD_LOGIC;
			q_n, q : out STD_LOGIC_VECTOR(7 downto 0);
			btn3 : in STD_LOGIC);
end component;


component bcd_converter is
    Port ( entrada : in  STD_LOGIC_VECTOR (7 downto 0);
           sum : out  STD_LOGIC_VECTOR (7 downto 0));
end component;


component rand_gen is
    Port ( clock, clock_2, btn3 : in  STD_LOGIC;
           q_n, q : out  STD_LOGIC_VECTOR (7 downto 0));
end component;


component comparator is
    Port ( a, b : in  STD_LOGIC_VECTOR (7 downto 0);
				btn1 : in STD_LOGIC;
           comp : out  STD_LOGIC);
end component;


component swf is
    Port ( switch : in  STD_LOGIC_VECTOR (7 downto 0);
           led : out  STD_LOGIC_VECTOR (7 downto 0));
end component;



begin


conversor : component bcd_converter
	port map(
		entrada => qr,
		sum => binario_aleatorio);


comparador : component comparator 
    Port map(
		a => binario_aleatorio,
		b => sw_s,
		btn1 => btn1,
		comp => confirmador);


switch_map : component swf 
	port map(
		switch => sw_s,
		led => led_s);


divisor : component div_f
	port map(
		clk_d => clock,
		reset => btn3,
		clk_1 => clk_1,
		clk_3 => clk_3,
		clk_250 => clk_250);


countdown : component countdowni
	port map(
		clock => clk_1,
		q_n => q_nc,
		q => qc,
		btn3 => btn3);
		

		
gerador : component rand_gen
	port map(
		clock => clk_250,
		clock_2 => clk_3,
		q_n => q_nr,
		q => qr,
		btn3 => btn3);
		


led <= led_s;
an <= an_s;
sw_s <= switch;
cx <= cx_s;


process(clk_250)
variable conta4 : integer := 1 ;
begin

	if rising_edge(clk_250) then
	
	
	if(conta4 = 1) then
		cx_s <= disp3;
		an_s <= "0111";
		conta4 := conta4 + 1;

		
	
	elsif(conta4 = 2) then 
		cx_s <= disp2;
		an_s <= "1011";
		conta4 := conta4 + 1;


	elsif(conta4 = 3) then
		cx_s <= disp1;
		an_s <= "1101";
		conta4 := conta4 + 1;

	
	elsif(conta4 = 4) then 
		cx_s <= disp0;
		an_s <= "1110";
		conta4 := 1;

end if;	
end if;
end process;



process(clk_250, qc, qr, chave, binario_aleatorio, sw_s, confirmador)
	begin
		
	if (btn1 = '1' ) then
		chave <= '0';
	end if;
		
		
	if(qc = "01000001") then
		disp0 <= "10001110"; 
		disp1 <= "10001110"; 
	else
	
	if(chave = '1') then
		case qc(3 downto 0) is
			when "0000" => disp0 <= "11000000"; --0
			when "0001" => disp0 <= "10010000"; --9
			when "0010" => disp0 <= "10000000"; --8
			when "0011" => disp0 <= "11111000"; --7
			when "0100" => disp0 <= "10000010"; --6
			when "0101" => disp0 <= "10010010"; --5
			when "0110" => disp0 <= "10011001"; --4
			when "0111" => disp0 <= "10110000"; --3
			when "1000" => disp0 <= "10100100"; --2
			when "1001" => disp0 <= "11111001"; --1
			when others => disp0 <= "11111111"; --APAGADO
		end case;
			
		case qc(7 downto 4) is
			when "0000" => disp1 <= "10110000"; --3
			when "0001" => disp1 <= "10100100"; --2
			when "0010" => disp1 <= "11111001"; --1
			when "0011" => disp1 <= "11000000"; --0
			when others => disp1 <= "11111111"; --APAGADO
		end case;
	elsif(chave = '0') then
		case confirmador is
			when '0' => disp0 <= "10001110"; 
							disp1 <= "10001110"; 
			when '1' => disp0 <= "10000010";
							disp1 <= "10000010";
			when others => disp1 <= "11111111";
								disp0 <= "11111111";
		end case;
	end if;
end if;


	case qr(3 downto 0) is
		when "0000" => disp2 <= "11000000"; --0
		when "0001" => disp2 <= "11111001"; --1
		when "0010" => disp2 <= "10100100"; --2
		when "0011" => disp2 <= "10110000"; --3
		when "0100" => disp2 <= "10011001"; --4
		when "0101" => disp2 <= "10010010"; --5
		when "0110" => disp2 <= "10000010"; --6
		when "0111" => disp2 <= "11111000"; --7
		when "1000" => disp2 <= "10000000"; --8
		when "1001" => disp2 <= "10010000"; --9
		when others => disp2 <= "11111111"; --APAGADO
	end case;
	
	case qr(7 downto 4) is
		when "0000" => disp3 <= "11000000"; --0
		when "0001" => disp3 <= "11111001"; --1
		when "0010" => disp3 <= "10100100"; --2
		when "0011" => disp3 <= "10110000"; --3
		when "0100" => disp3 <= "10011001"; --4
		when "0101" => disp3 <= "10010010"; --5
		when "0110" => disp3 <= "10000010"; --6
		when "0111" => disp3 <= "11111000"; --7
		when "1000" => disp3 <= "10000000"; --8
		when "1001" => disp3 <= "10010000"; --9
		when others => disp3 <= "11111111"; --APAGADO
	end case;
	
end process;



end Behavioral;

